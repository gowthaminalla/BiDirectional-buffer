* C:\Users\Gowthami\Desktop\ltspice\GPIO.asc
R1 N002 PUEN 10K
R2 PDEN 0 10K
XU1 PI Y PO NAND_2
V1 EN 0 PULSE(0 3.3 1m 1m 1m 0.5 1 5)
V2 N002 0 3.3
V3 N006 0 3.3
XU2 EN N003 INV_1
V4 A 0 PULSE(0 3.3 1m 1m 1m 0.5 1 5)
XU3 PDEN N010 INV_1
V7 N001 0 3.3
M1 N009 PUEN N001 N001 CMOSN NMOS l=12u w=3u
M3 N009 N010 0 0 CMOSP PMOS l=9u w=3u m=1
M4 N004 Y N003 N003 CMOSP PMOS l=9u w=3u m=1
M5 N007 A EN EN CMOSP PMOS l=9u w=3u m=1
M6 Y N007 EN EN CMOSP PMOS l=9u w=3u m=1
M7 A N004 0 0 CMOSN NMOS l=12u w=3u
M8 N004 Y 0 0 CMOSN NMOS l=12u w=3u
M9 N007 A 0 0 CMOSN NMOS l=12u w=3u
M10 Y N007 0 0 CMOSN NMOS l=12u w=3u
M2 A N004 N003 N003 CMOSP PMOS l=9u w=3u m=1
M11 PUEN N005 0 0 CMOSN NMOS l=12u w=3u
R3 N005 0 10K
M12 N006 N008 PDEN PDEN CMOSN NMOS l=12u w=3u
R4 N008 0 10K
.tran 0 8s 0s 0.1s
.include PMOS-180nm.lib
.include NMOS-180nm.lib
.lib DigitalLogic.lib
*control
.control
run
plot V(EN) 
plot V(Y)
plot V(A)
.endc
.end
