magic
tech scmos
timestamp 1594023687
<< metal1 >>
rect -63 70 -30 77
rect -63 69 -50 70
rect -84 59 -50 69
rect -15 61 -9 73
rect -164 26 -121 27
rect -164 20 -83 26
rect -159 19 -83 20
rect -159 -19 -150 19
rect -82 -1 -78 6
rect -159 -21 -149 -19
rect -159 -27 -135 -21
rect -82 -23 -73 -1
rect -101 -26 -73 -23
rect -63 -45 -50 59
rect -18 58 -9 61
rect -7 22 63 25
rect -11 17 63 22
rect -11 4 -5 17
rect 90 16 110 20
rect -15 -35 -10 -19
rect -15 -41 0 -35
rect -63 -50 -31 -45
rect -6 -46 0 -41
rect -51 -51 -31 -50
rect -1 -61 0 -46
<< m2contact >>
rect -83 19 -76 27
rect -78 -1 -73 6
rect -33 20 -26 26
rect -41 0 -34 6
<< metal2 >>
rect -76 21 -33 26
rect -73 0 -41 6
rect -73 -1 -36 0
use pmos  pmos_0
timestamp 1594014987
transform 1 0 -30 0 1 81
box -6 -9 24 29
use pmos  pmos_1
timestamp 1594014987
transform 1 0 -30 0 1 30
box -6 -9 24 29
use cmosinvereter  cmosinvereter_1
timestamp 1594009342
transform 1 0 -118 0 1 -26
box -18 -23 23 40
use nmos  nmos_0
timestamp 1594015197
transform 1 0 -17 0 1 -12
box -19 -11 12 17
use cmosinvereter  cmosinvereter_0
timestamp 1594009342
transform 1 0 80 0 1 17
box -18 -23 23 40
use nmos  nmos_1
timestamp 1594015197
transform 1 0 -13 0 1 -63
box -19 -11 12 17
<< labels >>
rlabel space -26 108 -26 108 5 vdd
rlabel space -12 -72 -12 -72 1 ground
rlabel space 76 54 76 54 1 vdd
rlabel space 83 -3 83 -3 1 ground
rlabel space -123 10 -122 10 1 vdd
rlabel space -116 -45 -116 -45 1 ground
rlabel metal1 -84 59 -84 69 1 vin
rlabel metal1 -164 20 -164 27 3 ven
rlabel metal1 110 16 110 20 7 vout
<< end >>
