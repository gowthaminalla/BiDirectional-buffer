* C:\Users\Gowthami\Desktop\ltspice\GPIO.asc
R1 N002 PUEN 10K
R2 PDEN 0 10K
V1 EN 0 PWL(0 1 1.9999 1 2 1 3.9999 1 4 1 5.9999 1 6 1 7.9999 1 8 1 9.9999 1 10 1 11.9999 1 12 1 13.9999 1 14 1 15.9999 1 16 1 17.9999 1 18 1 19.9999 1)
V4 A 0 PWL(0 0 1.9999 0 2 1.8 3.9999 1.8 4 1.8 5.9999 1.8 6 0 6.9999 0 7 1.8 7.9999 1.8 8 0 8.9999 0 9 1.8 9.9999 1.8 10 0 11.9999 0 12 1.8 13.9999 1.8 14 1.8 15.9999 1.8)
V7 N001 0 1.8
R3 N006 0 10K
R4 N008 0 10K
XX1 PDEN N010 inverter
XX3 PI Y PO nand
M5 Y N005 N003 N003 CMOSP l=180n w=900n m=1
M6 Y N005 0 0 CMOSN l=180n w=360n
M2 N005 N004 N003 N003 CMOSP l=180n w=900n m=1
M4 N005 N004 0 0 CMOSN l=180n w=360n
M7 PUEN N006 0 0 CMOSN l=180n w=360n
M8 N007 N008 PDEN PDEN CMOSN l=180n w=360n
M9 N009 PUEN N001 N001 CMOSN l=180n w=360n
M10 N009 N010 0 0 CMOSP l=180n w=900n m=1
V5 PI 0 PWL(0 0 0.9999 0 1 1.8 1.999 1.8 2 0 3.9999 0 4 1.8 5.9999 1.8 6 1.8 7.9999 1.8 8 0 9.9999 0 10 0 10.9999 0 11 1.8 11.9999 1.8 12 0 13.9999 0 14 1.8 15.9999 1.8)
XX2 A EN N004 tristate
V6 N003 0 1.8
V8 N002 0 PWL(0 0 0.9999 0 1 1.8 1.9999 1.8 2 0 2.9999 0 3 1.8 3.9999 1.8 4 0 4.9999 0 5 1.8 5.9999 1.8 6 1.8 7.9999 1.8 8 1.8 9.9999 1.8 10 1.8 11.9999 1.8 12 0 13.9999 0 14 0 15.9999 0)
V9 N007 0 PWL(0 0 0.9999 0 1 1.8 1.9999 1.8 2 0 2.9999 0 3 1.8 3.9999 1.8 4 0 4.9999 0 5 1.8 5.9999 1.8 6 1.8 7.9999 1.8 8 1.8 9.9999 1.8 10 0 11.9999 0 12 1.8 13.9999 1.8 14 1.8 15.9999 1.8)

* block symbol definitions
.subckt inverter I O
V1 N001 0 1.8
M1 O I N001 N001 CMOSP l=180n w=900n m=1
M2 O I 0 0 CMOSN l=180n w=360n
.include PMOS-180nm.lib
.include NMOS-180nm.lib
.ends inverter

.subckt nand A B O
V1 N001 0 1.8
M1 O A N001 N001 CMOSP l=180n w=900n m=1
M2 O B N001 N001 CMOSP l=180n w=900n m=1
M3 N002 B 0 0 CMOSN l=180n w=360n
M4 O A N002 0 CMOSN l=180n w=360n
.include NMOS-180nm.lib
.include PMOS-180nm.lib
.ends nand

.subckt tristate I EN O
V1 N001 0 1.8
M1 N003 EN N004 N004 CMOSP l=180n w=900n m=1
M2 N005 EN N001 N001 CMOSP l=180n w=900n m=1
M5 N004 I N001 N002 CMOSP l=180n w=900n m=1
M3 N003 N005 N006 N006 CMOSN l=180n w=360n
M4 N006 I 0 N007 CMOSN l=180n w=360n
M6 N005 EN 0 0 CMOSN l=180n w=360n
M7 O N003 N001 NC_01 CMOSP l=180n w=900n m=1
M8 O N003 0 0 CMOSN l=180n w=360n
.include PMOS-180nm.lib
.include NMOS-180nm.lib
.ends tristate
.tran 1 16s 0s 0.1s
.include PMOS-180nm.lib
.include NMOS-180nm.lib
* Tristate
* inverter
* NAND
*control
.control
run
plot V(EN) V(A)
plot V(PUEN) 
plot V(PDEN)
plot V(PO) V(PI) V(Y)
.endc
.end
