* C:\Users\Gowthami\Desktop\ltspice\GPIO with E=0.asc
R1 N002 PUEN 10K
V1 EN 0 PWL(0n 0 99.9999n 0)
V2 A 0 PWL(0n 0 49.9999n 0 50n 1.8 99.9999n 1.8)
V3 N001 0 1.8
R3 N006 0 10K
R4 N008 N007 10K
XX1 PDEN N010 inverter
XX2 PI Y PO nand
M1 Y N005 N003 N003 CMOSP l=180n w=900n m=1
M2 Y N005 0 0 CMOSN l=180n w=360n
M3 N005 N004 N003 N003 CMOSP l=180n w=900n m=1
M4 N005 N004 0 0 CMOSN l=180n w=360n
M5 PUEN N006 0 0 CMOSN l=180n w=360n
M6 N007 N008 PDEN PDEN CMOSN l=180n w=360n
M7 N009 PUEN N001 N001 CMOSN l=180n w=360n
M8 N009 N010 0 0 CMOSP l=180n w=900n m=1
V4 PI 0 PWL(0n 0 6.9999n 0 7n 1.8 13.9999n 1.8 14n 0 26.9999n 0 27n 1.8 39.9999n 1.8 40n 1.8 52.9999n 1.8 53n 0 65.9999n 0 66n 0 72.9999n 0 73n 1.8 79.9999n 1.8 80n 0 92.9999n 0 93n 1.8 102.9999n 1.8)
XX3 A EN N004 tristate
V5 N003 0 1.8
V6 N002 0 PWL(0n 0 6.9999n 0 7n 1.8 13.9999n 1.8 14n 0 20.9999n 0 21n 1.8 27.9999n 1.8 28n 0 34.9999n 0 35n 1.8 41.9999n 1.8 42n 1.8 54.9999n 1.8 55n 1.8 67.9999n 1.8 68n 1.8 80.9999n 1.8 81n 0 92.9999n 0 93n 0 99.9999n 0)
R2 PDEN 0 10K
V7 N007 0 PWL(0n 0 6.9999n 0 7n 1.8 13.9999n 1.8 14n 0 20.9999n 0 21n 1.8 27.9999n 1.8 28n 0 34.9999n 0 35n 1.8 41.9999n 1.8 42n 1.8 54.9999n 1.8 55n 1.8 67.9999n 1.8 68n 0 80.9999n 0 81n 1.8 92.9999n 1.8 93n 1.8 99.9999n 1.8)

* block symbol definitions
.subckt inverter I O
V1 N001 0 1.8
M1 O I N001 N001 CMOSP l=180n w=900n m=1
M2 O I 0 0 CMOSN l=180n w=360n
.include PMOS-180nm.lib
.include NMOS-180nm.lib
.ends inverter

.subckt nand A B O
V1 N001 0 1.8
M1 O A N001 N001 CMOSP l=180n w=900n m=1
M2 O B N001 N001 CMOSP l=180n w=900n m=1
M3 N002 B 0 0 CMOSN l=180n w=360n
M4 O A N002 0 CMOSN l=180n w=360n
.include NMOS-180nm.lib
.include PMOS-180nm.lib
.ends nand

.subckt tristate I EN O
V1 N001 0 1.8
M1 N003 EN N004 N004 CMOSP l=180n w=900n m=1
M2 N005 EN N001 N001 CMOSP l=180n w=900n m=1
M5 N004 I N001 N002 CMOSP l=180n w=900n m=1
M3 N003 N005 N006 N006 CMOSN l=180n w=360n
M4 N006 I 0 N007 CMOSN l=180n w=360n
M6 N005 EN 0 0 CMOSN l=180n w=360n
M7 O N003 N001 N001 CMOSP l=180n w=900n m=1
M8 O N003 0 0 CMOSN l=180n w=360n
.include PMOS-180nm.lib
.include NMOS-180nm.lib
.ends tristate
.tran 1 100n 0
.include PMOS-180nm.lib
.include NMOS-180nm.lib
* Tristate
* inverter
* NAND
*control
.control
run
plot V(EN)  V(A) V(Y)
.endc
.end

