* SPICE3 file created from bidir.ext - technology: scmos

.option scale=0.1u

M1000 m1_16_34# porta en cmosinvereter_0/w_n14_4# pfet w=7 l=3
+  ad=77 pd=36 as=537 ps=356
M1001 m1_16_34# porta cmosinvereter_0/a_n6_n8# en nfet w=5 l=3
+  ad=65 pd=36 as=77 ps=60
M1002 portb m1_16_34# en cmosinvereter_1/w_n14_4# pfet w=7 l=3
+  ad=154 pd=72 as=0 ps=0
M1003 portb m1_16_34# cmosinvereter_1/a_n6_n8# en nfet w=5 l=3
+  ad=130 pd=72 as=77 ps=60
M1004 m1_19_n46# porta en cmosinvereter_2/w_n14_4# pfet w=7 l=3
+  ad=77 pd=36 as=0 ps=0
M1005 m1_19_n46# porta cmosinvereter_2/a_n6_n8# en nfet w=5 l=3
+  ad=65 pd=36 as=77 ps=60
M1006 portb m1_19_n46# en cmosinvereter_3/w_n14_4# pfet w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1007 portb m1_19_n46# cmosinvereter_3/a_n6_n8# en nfet w=5 l=3
+  ad=0 pd=0 as=77 ps=60
M1008 en en en cmosinvereter_4/w_n14_4# pfet w=7 l=3
+  ad=0 pd=0 as=0 ps=0
M1009 en en cmosinvereter_4/a_n6_n8# en nfet w=5 l=3
+  ad=65 pd=36 as=77 ps=60
