magic
tech scmos
timestamp 1594012772
<< metal1 >>
rect -113 77 59 82
rect -113 75 47 77
rect -112 60 -104 75
rect -42 74 -10 75
rect -131 49 -104 60
rect -112 19 -104 49
rect -28 34 -19 38
rect 38 37 46 40
rect 16 34 46 37
rect 79 36 105 40
rect -112 15 -94 19
rect -59 14 -34 17
rect -46 7 -34 14
rect -46 0 -40 7
rect -28 -32 -20 34
rect 100 16 104 36
rect 100 6 112 16
rect 4 3 66 6
rect -2 -5 4 0
rect 62 -1 66 3
rect -43 -42 -20 -32
rect 100 -36 104 6
rect 48 -42 54 -38
rect 96 -39 104 -36
rect 85 -42 104 -39
rect -28 -46 -16 -42
rect 48 -43 58 -42
rect 19 -46 58 -43
rect -28 -47 -20 -46
<< m2contact >>
rect -40 0 -34 7
rect -2 0 4 6
<< metal2 >>
rect -40 7 4 8
rect -34 6 4 7
rect -34 0 -2 6
use cmosinvereter  cmosinvereter_4
timestamp 1594012772
transform 1 0 -76 0 1 16
box -18 -23 23 40
use cmosinvereter  cmosinvereter_0
timestamp 1594012772
transform 1 0 -1 0 1 35
box -18 -23 23 40
use cmosinvereter  cmosinvereter_1
timestamp 1594012772
transform 1 0 62 0 1 37
box -18 -23 23 40
use cmosinvereter  cmosinvereter_2
timestamp 1594012772
transform 1 0 2 0 1 -45
box -18 -23 23 40
use cmosinvereter  cmosinvereter_3
timestamp 1594012772
transform 1 0 69 0 1 -41
box -18 -23 23 40
<< labels >>
rlabel metal1 -131 49 -131 60 3 en
rlabel metal1 112 6 112 16 7 portb
rlabel metal1 -43 -42 -43 -32 1 porta
rlabel space 4 -64 4 -64 1 gnd
rlabel space 72 -60 72 -60 1 gnd
rlabel space 64 16 64 16 1 gnd
rlabel space 2 16 2 16 1 gnd
<< end >>
