magic
tech scmos
timestamp 1594009342
<< nwell >>
rect -14 4 23 29
<< ntransistor >>
rect 2 -8 5 -3
<< ptransistor >>
rect 2 10 5 17
<< ndiffusion >>
rect -6 -4 2 -3
rect -6 -8 -5 -4
rect 0 -8 2 -4
rect 5 -7 11 -3
rect 15 -7 18 -3
rect 5 -8 18 -7
<< pdiffusion >>
rect -2 14 2 17
rect -6 10 2 14
rect 5 16 16 17
rect 5 12 10 16
rect 14 12 16 16
rect 5 10 16 12
<< ndcontact >>
rect -5 -9 0 -4
rect 11 -7 15 -3
<< pdcontact >>
rect -6 14 -2 18
rect 10 12 14 16
<< psubstratepcontact >>
rect -12 34 -8 38
rect 1 34 5 38
<< nsubstratencontact >>
rect -5 -22 -1 -18
rect 6 -22 10 -18
<< polysilicon >>
rect 2 17 5 23
rect 2 2 5 10
rect -7 -1 5 2
rect 2 -3 5 -1
rect 2 -10 5 -8
<< polycontact >>
rect -11 -1 -7 3
<< metal1 >>
rect -15 38 10 40
rect -15 34 -12 38
rect -8 34 1 38
rect 5 34 10 38
rect -15 29 10 34
rect -14 24 10 29
rect -14 18 1 24
rect -14 14 -6 18
rect -2 14 1 18
rect 14 12 17 16
rect -18 -1 -11 3
rect 10 -3 17 12
rect -6 -9 -5 -6
rect 10 -7 11 -3
rect 15 -7 17 -3
rect -6 -13 0 -9
rect -6 -18 13 -13
rect -6 -22 -5 -18
rect -1 -22 6 -18
rect 10 -22 13 -18
rect -6 -23 13 -22
<< end >>
