* C:\Users\Gowthami\Desktop\ltspice\GPIO.asc
R1 N002 PUEN 10K
R2 PDEN 0 10K
XU1 PI Y PO NAND_2
V1 EN 0 PULSE(0 3.3 10m 1n 1n 10m 20m 10)
V2 N002 0 3.3
V3 N006 0 3.3
XU2 EN N003 INV_1
V4 A 0 PULSE(0 3.3 10m 1n 1n 10m 20m 10)
XU3 PDEN N010 INV_1
V7 N001 0 3.3
M1 N009 PUEN N001 N001 CMOSN l=180n w=360n
M3 N009 N010 0 0 CMOSP l=180n w=900n m=1
M4 N004 Y N003 N003 CMOSP l=180n w=900n m=1
M5 N007 A EN EN CMOSP l=180n w=900n m=1
M6 Y N007 EN EN CMOSP l=180n w=900n m=1
M7 A N004 0 0 CMOSN l=180n w=360n
M8 N004 Y 0 0 CMOSN l=180n w=360n
M9 N007 A 0 0 CMOSN l=180n w=360n
M10 Y N007 0 0 CMOSN l=180n w=360n
M2 A N004 N003 N003 CMOSP l=180n w=900n m=1
M11 PUEN N005 0 0 CMOSN l=180n w=360n
R3 N005 0 10K
M12 N006 N008 PDEN PDEN CMOSN l=180n w=360n
R4 N008 0 10K
.tran 0 8s 0s 0.1s
.include PMOS-180nm.lib
.include NMOS-180nm.lib
.lib DigitalLogic.lib
*control
.control
run
plot V(EN) 
plot V(Y)
plot V(A)
.endc
.end
