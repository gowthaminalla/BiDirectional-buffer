magic
tech scmos
timestamp 1593856735
<< nwell >>
rect -8 4 15 29
<< ntransistor >>
rect 2 -8 5 -3
<< ptransistor >>
rect 2 10 5 17
<< ndiffusion >>
rect -6 -8 2 -3
rect 5 -8 13 -3
<< pdiffusion >>
rect -2 10 2 17
rect 5 10 9 17
<< polysilicon >>
rect 2 17 5 23
rect 2 -3 5 10
rect 2 -10 5 -8
<< metal1 >>
rect -8 24 10 29
rect -8 18 1 24
rect -2 14 1 18
rect -6 -13 0 -6
rect -6 -18 13 -13
<< end >>
